`ifndef PKT_DEC_SV
`define PKT_DEC_SV

class pkt_dec;
	
	parameter DATA_WD = 8;
	
endclass

`endif